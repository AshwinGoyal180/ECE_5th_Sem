library ieee;
use ieee.std_logic_1164.all;

entity sub_tb is
end sub_tb;

architecture ADDER of sub_tb is
    component fullsubtractor is
        port (
            A  : in  std_logic;
            B  : in  std_logic;
            C : in  std_logic;
            D  : out std_logic;
            BO : out std_logic);
    end component;
    signal input  : std_logic_vector(2 downto 0);
    signal output : std_logic_vector(1 downto 0);
begin
    uut: fullsubtractor port map (
        A => input(2),
        B => input(1),
        C => input(0),
        D => output(0),
        BO => output(1)
    );

    stim_proc: process
    begin
        input <= "000"; wait for 10 ns; assert output = "00" report "0+0+0 failed";
        input <= "001"; wait for 10 ns; assert output = "11" report "0+0+1 failed";
        input <= "010"; wait for 10 ns; assert output = "11" report "0+1+0 failed";
        input <= "011"; wait for 10 ns; assert output = "10" report "0+1+1 failed";
        input <= "100"; wait for 10 ns; assert output = "01" report "1+0+0 failed";
        input <= "101"; wait for 10 ns; assert output = "00" report "1+0+1 failed";
        input <= "110"; wait for 10 ns; assert output = "00" report "1+1+0 failed";
        input <= "111"; wait for 10 ns; assert output = "11" report "1+1+1 failed";
        report "Full subtractor testbench finished";
        wait;
    end process;
end;
